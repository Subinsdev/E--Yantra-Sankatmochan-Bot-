module color_sense(
						input clk,
						input c_clk,
						output [2:0]color,
						output s2,
						output s3
);
	
	parameter IDLE = 3'b000;
	parameter RED_START = 3'b001;
	parameter RED_READ = 3'b010;
	parameter GREEN_START = 3'b011;
	parameter GREEN_READ = 3'b100;
	parameter BLUE_START = 3'b101;
	parameter BLUE_READ = 3'b110;
	
	// set the thresholds here
	// To test the program is correct or not please simulate waveform6.vwf with these thresholds and the specified parameters
	parameter R_THRESH_HIGH = 120;
	parameter R_THRESH_LOW = 25;
	parameter G_THRESH_HIGH = 120;
	parameter G_THRESH_LOW = 25;
	parameter B_THRESH_HIGH = 120;
	parameter B_THRESH_LOW = 25;
	
	reg [8:0]counter;
	reg [8:0]c_counter;
	reg [2:0]r_state = IDLE;
	reg [1:0]out_color = 0;
	reg out_s2 = 1;
	reg out_s3 = 0;
	
	always @(posedge clk)
		begin
			case(r_state)
				IDLE :
					begin
						out_color <= 0;
						out_s2 <= 1;
						out_s3 <= 0;
						r_state <= RED_START;
					end
				RED_START :
					begin
						out_s2 <= 0;
						out_s3 <= 0;
						counter <= 0;
						
						r_state <= RED_READ;
					end
				RED_READ :
					begin
						if(counter < 300)
						begin
							counter <= counter + 1'b1;
							r_state <= RED_READ;
						end
						else
						begin
							r_state <= GREEN_START;
							if(c_counter < R_THRESH_HIGH && c_counter > R_THRESH_LOW)
								out_color <= 1;
						end
						
					end
				GREEN_START :
					begin
						out_s2 <= 1;
						out_s3 <= 1;
						counter <= 0;
						r_state <= GREEN_READ;
					end
				GREEN_READ :
					begin
						if(counter < 300)
						begin
							counter <= counter + 1'b1;
							r_state <= GREEN_READ;
						end
						else
						begin
							r_state <= BLUE_START;
							if(c_counter < G_THRESH_HIGH && c_counter > G_THRESH_LOW)
								out_color <= 2;
						end
						
					end
				BLUE_START :
					begin
						out_s2 <= 0;
						out_s3 <= 1;
						counter <= 0;
						r_state <= BLUE_READ;
					end
				BLUE_READ :
					begin
						if(counter < 300)
						begin
							counter <= counter + 1'b1;
							r_state <= BLUE_READ;
						end
						else
						begin
							r_state <= IDLE;
							if(c_counter < B_THRESH_HIGH && c_counter > B_THRESH_LOW)
								out_color <= 3;
						end
						
					end
				
			endcase
			
		end
	
	always@(posedge c_clk)
		begin
			c_counter <= c_counter + 1'b1;
			if(counter == 0)
			begin
				$display("max c_counter: 0x%0h", c_counter);
				c_counter <= 0;
			end
		end
								
	assign color = out_color;
	assign s2 = out_s2;
	assign s3 = out_s3;
	
endmodule
	